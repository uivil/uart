module debouncer (input in, output out);

assign out = in;

endmodule
